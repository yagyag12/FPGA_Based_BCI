/************************************************************/
//           W I N D O W I N G   M O D U L E                //
//                                                          //
//  Desc: Does Hamming windowing for preventing leakage     //
/************************************************************/
`timescale 1ns / 1ps

module windowing_module #(
    parameter EPOCH_LENGTH = 256
)(
    input                       clk,
    input                       rst,
    input                       en,
    input  logic signed [31:0]  signal_in,
    output logic signed [31:0]  windowed_signal,
    output logic                o_window_done,
    output logic                o_window_valid
    );

/***********************  SIGNALS  **************************/

// Window Coefficients 
logic signed [15:0] window_coeffs [0:255] = '{
    1311, 1313, 1320, 1331, 1347, 1368, 1393, 1423, 1457, 1495, 1538, 1586, 1638, 1694, 1755, 1820,
    1889, 1962, 2040, 2122, 2207, 2297, 2391, 2489, 2591, 2696, 2805, 2918, 3034, 3154, 3278, 3405,
    3535, 3668, 3804, 3944, 4086, 4232, 4380, 4531, 4684, 4840, 4999, 5160, 5323, 5488, 5655, 5824,
    5995, 6168, 6343, 6518, 6696, 6874, 7054, 7235, 7417, 7600, 7783, 7967, 8152, 8337, 8522, 8708,
    8894, 9079, 9265, 9450, 9635, 9820, 10003, 10187, 10369, 10550, 10731, 10910, 11088, 11264, 11440, 11613,
    11785, 11955, 12123, 12290, 12454, 12616, 12775, 12933, 13087, 13240, 13389, 13536, 13680, 13821, 13959, 14094,
    14226, 14354, 14479, 14601, 14719, 14834, 14945, 15052, 15155, 15255, 15351, 15443, 15531, 15614, 15694, 15770,
    15841, 15908, 15971, 16029, 16083, 16133, 16178, 16219, 16256, 16288, 16315, 16338, 16356, 16370, 16379, 16383,
    16383, 16379, 16370, 16356, 16338, 16315, 16288, 16256, 16219, 16178, 16133, 16083, 16029, 15971, 15908, 15841,
    15770, 15694, 15614, 15531, 15443, 15351, 15255, 15155, 15052, 14945, 14834, 14719, 14601, 14479, 14354, 14226,
    14094, 13959, 13821, 13680, 13536, 13389, 13240, 13087, 12933, 12775, 12616, 12454, 12290, 12123, 11955, 11785,
    11613, 11440, 11264, 11088, 10910, 10731, 10550, 10369, 10187, 10003, 9820, 9635, 9450, 9265, 9079, 8894,
    8708, 8522, 8337, 8152, 7967, 7783, 7600, 7417, 7235, 7054, 6874, 6696, 6518, 6343, 6168, 5995,
    5824, 5655, 5488, 5323, 5160, 4999, 4840, 4684, 4531, 4380, 4232, 4086, 3944, 3804, 3668, 3535,
    3405, 3278, 3154, 3034, 2918, 2805, 2696, 2591, 2489, 2391, 2297, 2207, 2122, 2040, 1962, 1889,
    1820, 1755, 1694, 1638, 1586, 1538, 1495, 1457, 1423, 1393, 1368, 1347, 1331, 1320, 1313, 1311
};

logic        [$clog2(EPOCH_LENGTH):0] window_idx;
logic signed [63:0]                   windowed_signal_acc;


/**********************  WINDOWING  *************************/

always_ff @(posedge clk or posedge rst) begin
    if (rst) begin
        windowed_signal_acc <= 0;
        o_window_done       <= 0;
        o_window_valid      <= 0;
        window_idx          <= 0;
    end 
    else if (en) begin
        if (window_idx < EPOCH_LENGTH) begin
            windowed_signal_acc <= signal_in * window_coeffs[window_idx];
            o_window_valid      <= 1;
            window_idx          <= window_idx + 1;
            o_window_done       <= 0;
        end 
        else begin
            windowed_signal_acc <= 0;
            o_window_valid      <= 0;
            o_window_done       <= 1;
            window_idx          <= 0;
        end
    end 
    else begin
        o_window_done   <= 0;
        o_window_valid  <= 0; 
    end
end

assign windowed_signal = {windowed_signal_acc[63], windowed_signal_acc[59:28]};

endmodule
